-- SP next move on the FPGA
--
-- entity name: g29_sp_next_move
--
-- Version 1.1
-- Author: Stepan Salenikovich, Ayman Zakir
-- Date: 25.11.2011

-- INSTRUCTIONS (key mappings):
-- SW[9 - 7] - input GRA row
-- SW[6 - 4] - input GRA col
-- SW[1,0] - input GRA[1,0]
-- KEY3 - write to GRA
-- KEY0 - reset
-- LEDR[9 - 4, 1, 0] - light up when corresponding switches are high
-- HEX3 - selected GRA row
-- HEX2 - selected GRA col
-- HEX[1,0] - contents of selected GRA[1,0]

library ieee; -- allows use of the std_logic_vector type
use ieee.std_logic_1164.all;

entity g29_FPGA_sp_next_move is
	port(
		-- NM, ASPMC: in std_logic;
		-- cyclone II board I/O
		SW_row, SW_col: in natural range 0 to 7;
		SW_gra_value: in std_logic_vector(0 to 1);
		KEY_write, KEY_reset: in std_logic; -- push to write
		LEDR_row, LEDR_col: out natural range 0 to 7; -- LEDs light up when value high
		LEDR_gra_value: out std_logic_vector(0 to 1);
		--
		clk: in std_logic;
		-- rst: in std_logic;
		mc_count: out natural range 0 to 16;
		SPMC: out std_logic;
		-- 7 seg LED displays
		HEX0: out std_logic_vector(6 downto 0);
		HEX1: out std_logic_vector(6 downto 0);
		HEX2: out std_logic_vector(6 downto 0);
		HEX3: out std_logic_vector(6 downto 0)
	);
end g29_FPGA_sp_next_move;

architecture concurrent of g29_FPGA_sp_next_move is

	-- Generated by Quartus II Version 9.0 (Build Build 235 06/17/2009)
	-- Created on Fri Nov 25 15:09:18 2011

	COMPONENT g29_sp_player
		PORT
		(
			NM				:	 IN STD_LOGIC;
			ASPMC			:	 IN STD_LOGIC;
			gra_read		:	 IN STD_LOGIC_VECTOR(0 TO 1);
			write_enable	:	 OUT STD_LOGIC;
			gra_row			:	 OUT NATURAL RANGE 0 TO 7;
			gra_col			:	 OUT NATURAL RANGE 0 TO 7;
			gra_write		:	 OUT STD_LOGIC_VECTOR(0 TO 1);
			SW_row			:	 IN NATURAL RANGE 0 TO 7;
			SW_col			:	 IN NATURAL RANGE 0 TO 7;
			SW_gra_value	:	 IN STD_LOGIC_VECTOR(0 TO 1);
			KEY_write		:	 IN STD_LOGIC;
			clk				:	 IN STD_LOGIC;
			rst				:	 IN STD_LOGIC;
			mc_count		:	 OUT NATURAL RANGE 0 TO 31;
			SPMC			:	 OUT STD_LOGIC
		);
	END COMPONENT;
	
	-- Generated by Quartus II Version 9.0 (Build Build 235 06/17/2009)
	-- Created on Fri Nov 25 15:18:47 2011

	COMPONENT g29_gra_arr
		PORT
		(
			row_in			:	 IN NATURAL RANGE 0 TO 7;
			col_in			:	 IN NATURAL RANGE 0 TO 7;
			gra_in			:	 IN STD_LOGIC_VECTOR(0 TO 1);
			write_enable	:	 IN STD_LOGIC;
			clk				:	 IN STD_LOGIC;
			rst				:	 IN STD_LOGIC;
			gra_out			:	 OUT STD_LOGIC_VECTOR(0 TO 1)
		);
	END COMPONENT;

-- Generated by Quartus II Version 9.0 (Build Build 235 06/17/2009)
-- Created on Fri Nov 25 16:45:33 2011

COMPONENT g29_7_segment_decoder
	PORT
	(
		clk					:	 IN STD_LOGIC;
		number				:	 IN NATURAL RANGE 0 TO 7;
		seven_seg_display	:	 OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;
	-- end generated code
	
	signal row, col : natural range 0 to 7;
	signal gra_read, gra_write : std_logic_vector(0 to 1);
	signal write_enable : std_logic;
	signal h0, h1 : natural range 0 to 7;
	
begin
	
	player : g29_sp_player port map (	'0',
										'1',
										gra_read,
										write_enable,
										row,
										col,
										gra_write,
										SW_row,
										SW_col,
										SW_gra_value,
										KEY_write,
										clk,
										KEY_reset,
										mc_count,
										SPMC	);
										
	gra : g29_gra_arr port map (	row,
									col,
									gra_write,
									write_enable,
									clk,
									KEY_reset,
									gra_read	);
									
	h0 <= 1 when gra_read(1) = '1' else 0;
	h1 <= 1 when gra_read(0) = '1' else 0;
	
	diplay3 : g29_7_segment_decoder port map (	clk,
												SW_row,
												HEX3	);
												
	diplay2 : g29_7_segment_decoder port map (	clk,
												SW_col,
												HEX2	);
												
	diplay1 : g29_7_segment_decoder port map (	clk,
												h0,
												HEX1	);
												
	diplay0 : g29_7_segment_decoder port map (	clk,
												h1,
												HEX0	);
												
	LEDR_row <= SW_row;
	LEDR_col <= SW_col;
	LEDR_gra_value <= SW_gra_value;
	
end concurrent;